LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FF_JK IS
PORT( D, Clk, En : IN STD_LOGIC;
	Q : OUT STD_LOGIC );
END FF_JK;

ARCHITECTURE JK OF FF_JK IS
BEGIN
	PROCESS(CLK)
	BEGIN
		IF En = '0' THEN
			NULL;
		ELSIF RISING_EDGE(CLK) THEN
			Q <= D;
		END IF;
	END PROCESS;
END JK;