-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Fri Sep 16 17:58:23 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY L0902 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        W : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC;
        Qn : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        Qn1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END L0902;

ARCHITECTURE BEHAVIOR OF L0902 IS
    TYPE type_fstate IS (A,B,C,D);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,W)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            z <= '0';
            Qn <= "00";
            Qn1 <= "00";
        ELSE
            z <= '0';
            Qn <= "00";
            Qn1 <= "00";
            CASE fstate IS
                WHEN A =>
                    IF (NOT((W = '1'))) THEN
                        reg_fstate <= A;
                    ELSIF ((W = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    IF (NOT((W = '1'))) THEN
                        Qn1 <= "00";
                    ELSIF ((W = '1')) THEN
                        Qn1 <= "01";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Qn1 <= "00";
                    END IF;

                    Qn <= "00";

                    z <= '0';
                WHEN B =>
                    IF (NOT((W = '1'))) THEN
                        reg_fstate <= A;
                    ELSIF ((W = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;

                    IF (NOT((W = '1'))) THEN
                        Qn1 <= "00";
                    ELSIF ((W = '1')) THEN
                        Qn1 <= "10";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Qn1 <= "00";
                    END IF;

                    Qn <= "01";

                    z <= '0';
                WHEN C =>
                    IF (NOT((W = '1'))) THEN
                        reg_fstate <= D;
                    ELSIF ((W = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    IF ((W = '1')) THEN
                        Qn1 <= "10";
                    ELSIF (NOT((W = '1'))) THEN
                        Qn1 <= "11";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Qn1 <= "00";
                    END IF;

                    Qn <= "10";

                    z <= '1';
                WHEN D =>
                    IF (NOT((W = '1'))) THEN
                        reg_fstate <= A;
                    ELSIF ((W = '1')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D;
                    END IF;

                    IF (NOT((W = '1'))) THEN
                        Qn1 <= "00";
                    ELSIF ((W = '1')) THEN
                        Qn1 <= "11";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Qn1 <= "00";
                    END IF;

                    Qn <= "11";

                    z <= '1';
                WHEN OTHERS => 
                    z <= 'X';
                    Qn <= "XX";
                    Qn1 <= "XX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
